----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 19.02.2016 19:26:44
-- Design Name: 
-- Module Name: simpleDualPortMemory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.MAIN_DEFINITIONS.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DualPortMemory is
    Port ( 
	        CLK    : in   STD_LOGIC;
	        Addr_A : in   STD_LOGIC_VECTOR (PC_WIDTH-1 downto 0);
	        DO_A   : out  STD_LOGIC_VECTOR (WORD_WIDTH-1 downto 0);
	        WE_B   : in   STD_LOGIC;
	        Addr_B : in   STD_LOGIC_VECTOR (PC_WIDTH-1 downto 0);
	        DI_B   : in   STD_LOGIC_VECTOR (WORD_WIDTH-1 downto 0);
	        DO_B   : out  STD_LOGIC_VECTOR (WORD_WIDTH-1 downto 0)
			  );
end DualPortMemory;

architecture Behavioral of DualPortMemory is

-- declare a matrix of bits... the memory
type MEM_TYPE is array (0 to (2**(PC_WIDTH-2))-1) of std_logic_vector(WORD_WIDTH-1 downto 0);

constant InitValue0 : MEM_TYPE := (
			0 => "001000" & "00001" & "00000" & "11111" & "11111111111", -- ADDI    R1,R0,#-1      R1 <- (0)  + (-1)     = -1 (C=0)
        1 => "001001" & "00010" & "00000" & "00010" & "11111111101", -- RSUBI   R2,R0,#2		  R2 <- (0) - (-1)     = -2 (C=0)
        2 => "000111" & "00011" & "00000" & "00100" & "00000000000", -- RSUBKC  R3,R0,R4       R3 <- (-2) + /(0) +C  = -3
        3 => "000011" & "00100" & "00000" & "00001" & "00000000000", -- RSUBC   R4,R0,R1       R4 <- (-1) + /(0) +C  = -2 (C=1)
--	    0 => "001000" & "00001" & "00000" & "11111" & "11111111111", -- ADDI    R1,R0,#-1      R1 <- (0)  + (-1)     = -1 (C=0)
--        1 => "001001" & "00010" & "00001" & "11111" & "11111111101", -- RSUBI   R2,R1,#-3      R2 <- (-3) - (-1)     = -2 (C=0)
--        2 => "000111" & "00011" & "00000" & "00010" & "00000000000", -- RSUBKC  R3,R0,R2       R3 <- (-2) + /(0) +C  = -3
--        3 => "000011" & "00100" & "00000" & "00001" & "00000000000", -- RSUBC   R4,R0,R1       R4 <- (-1) + /(0) +C  = -2 (C=1)
        4 => "000010" & "00100" & "00100" & "00011" & "00000000000", -- ADDC    R4,R4,R3       R4 <- (-2) + (-3) +C  = -4 (C=1)
        5 => "000000" & "00101" & "00100" & "00001" & "00000000000", -- ADD     R5,R4,R1       R5 <- (-4) + (-1)     = -5 (C=1)
        6 => "000011" & "00110" & "00101" & "00001" & "00000000000", -- RSUBC   R6,R5,R1       R6 <- (-1) + /(-5)+C  = +4 (C=0)
        7 => "000001" & "00110" & "00110" & "00010" & "00000000000", -- RSUB    R6,R6,R2       R6 <- (-2) - (+4)     = -6 (C=1)
        8 => "001110" & "00111" & "00000" & "11111" & "11111111001", -- ADDIKC  R7,R0,#-7      R7 <- (0)  + (-7) +C  = -6
        9 => "001010" & "01000" & "00111" & "11111" & "11111111110", -- ADDIC   R8,R7,#-2      R8 <- (-6) + (-2) +C  = -7 (C=1)
        10 => "000101" & "01001" & "01000" & "00000" & "00000000001", -- CMP     R9,R8,R0       R9 <- (0)  - (-7)     = sign positive
        11 => "000101" & "01001" & "01000" & "00000" & "00000000011", -- CMPU    R9,R8,R0       R5 <- (0)  - (-7)     = sign negative
        12 => "101110" & "00000" & "00000" & "00000" & "00000100000", -- BRI     =>20           PC <-- PC + 8*4
        ---------------------------------------------------------------------------------------------------------------------------
        20 => "101100" & "00000" & "00000" & "01111" & "11111111111", -- IMM     x7FFF          IMM<-- x7FFF
        21 => "101000" & "00001" & "00000" & "11111" & "11111111111", -- ORI     R1,R0,#-1      R1 <-- x7FFFFFFF (sign positive)
        22 => "101100" & "00000" & "00000" & "10000" & "00000000000", -- IMM     x8000          IMM<-- x8000 
        23 => "001000" & "00010" & "00000" & "00000" & "00000000000", -- ADDI    R2,R0,#0       R2 <-- x80000000 (sign negative)
        24 => "101100" & "00000" & "00000" & "10000" & "00000000000", -- IMM     x8000          IMM<-- x8000 
        25 => "101011" & "00011" & "00001" & "11111" & "11111111111", -- ANDNI   R3,R1,#xFFFF   R3 <-- x7FFF0000 (sign positive)
        26 => "101100" & "00000" & "00000" & "01111" & "11111111111", -- IMM     x8000          IMM<-- x7FFF 
        27 => "101010" & "00100" & "00011" & "00000" & "00000000000", -- XORI    R4,R3,#xFFFF   R4 <-- x00000000 (sign positive)
        28 => "101111" & "00000" & "00100" & "00000" & "00000001000", -- BEQI    =>30           PC <-- PC + 2*4
        29 => "101110" & "00000" & "00000" & "11111" & "11111011100", -- BRI     =>20           PC <-- PC - 9*4
        ---------------------------------------------------------------------------------------------------------------------------
        30 => "001000" & "00001" & "00000" & "11111" & "11111111110", -- ADDI    R1,R0,#-2      R1 <-- -2
        31 => "010000" & "00010" & "00001" & "00001" & "00000000000", -- MUL     R2,R1,R1       R2 <-- +4
        32 => "010000" & "00011" & "00001" & "00001" & "00000000001", -- MULH    R3,R1,R1       R3 <-- 0
        33 => "010000" & "00100" & "00001" & "00001" & "00000000011", -- MULHU   R4,R1,R1       R4 <-- -4
        34 => "010000" & "00101" & "00010" & "00001" & "00000000010", -- MULHSU  R5,R2,R4       R5 <-- +3
        35 => "101110" & "00010" & "01100" & "00000" & "00010010100", -- BRALI   R2,==>37       R2 <-- 140, PC <-- 37x4
        36 => "100110" & "00000" & "01000" & "00000" & "00000000000", -- BRA     R0             PC <-- 0
        37 => "100111" & "00100" & "00001" & "00000" & "00000000000", -- BGT     R1,R0          PC <-- PC + 4
        38 => "100111" & "00101" & "00001" & "00000" & "00000000000", -- BGE     R1,R0          PC <-- PC + 4
        39 => "100111" & "00011" & "00010" & "00000" & "00000000000", -- BLE     R2,R0          PC <-- PC + 4
        ---------------------------------------------------------------------------------------------------------------------------
        40 => "001000" & "00001" & "00000" & "11111" & "11100000001", -- ADDI    R1,R0,#xFF01   R1 <-- 0xFFFFFF01
        41 => "100100" & "00010" & "00001" & "00000" & "00001100001", -- SEXT16  R2,R1          R2 <-- 0xFFFFFF01
        42 => "100100" & "00011" & "00010" & "00000" & "00001100000", -- SEXT8   R3,R2          R3 <-- 0x00000001
        43 => "100100" & "00100" & "00010" & "00000" & "00001000001", -- SRL     R4,R2          R4 <-- 0x7FFFFF80 (C=1)
        44 => "100100" & "00101" & "00010" & "00000" & "00001000001", -- SRL     R5,R2          R5 <-- 0x7FFFFF80 (C=1)
        45 => "100100" & "00110" & "00100" & "00000" & "00000100001", -- SRC     R6,R4          R6 <-- 0xBFFFFFC0 (C=0)
        46 => "100100" & "00111" & "00110" & "00000" & "00000100001", -- SRC     R7,R6          R7 <-- 0x5FFFFFE0 (C=0)
        47 => "100100" & "01000" & "00110" & "00000" & "00000000001", -- SRA     R8,R6          R8 <-- 0xDFFFFFE0 (C=0)
        48 => "100100" & "01001" & "00111" & "00000" & "00000000001", -- SRA     R9,R7          R9 <-- 0x2FFFFFF0 (C=0)
        49 => "000000" & "00000" & "00001" & "00001" & "00000000000", -- ADD     R0,R1,R1       R0 <-- 0 (NOP)
        ---------------------------------------------------------------------------------------------------------------------------
        50 => "101100" & "00000" & "00000" & "01111" & "11111111111", -- IMM     x7FFF          IMM<-- x7FFF
        51 => "101000" & "00001" & "00000" & "11110" & "00000001111", -- ORI     R1,R0,#xF00F   R1 <-- x7FFFF00F
        52 => "101000" & "00010" & "00000" & "00000" & "00110010000", -- ORI     R2,R0,#400     R2 <-- 400
        53 => "110100" & "00001" & "00010" & "00000" & "00000000000", -- SB      (R0+R2),R1     M[400] <-- 0x0F
        54 => "111100" & "00001" & "00010" & "00000" & "00000000101", -- SBI     5(R2),R1       M[405] <-- 0x0F
        55 => "111100" & "00001" & "00010" & "00000" & "00000001010", -- SBI     10(R2),R1      M[410] <-- 0x0F
        56 => "111100" & "00001" & "00010" & "00000" & "00000001111", -- SBI     15(R2),R1      M[415] <-- 0x0F
        57 => "111101" & "00001" & "00010" & "00000" & "00000000010", -- SHI     2(R2),R1       M[402] <-- 0xF00F
        58 => "111110" & "00001" & "00010" & "00000" & "00000010000", -- SWI     16(R2),R1      M[416] <-- 0x7FFFF00F
        59 => "111001" & "00011" & "00010" & "00000" & "00000000100", -- LHUI    R3,4(R2)       R3 <-- 0x00000F00
        60 => "111001" & "00100" & "00010" & "00000" & "00000001010", -- LHUI    R4,10(R2)      R4 <-- 0x0000000F
        61 => "110010" & "00101" & "00010" & "00000" & "00000000000", -- LW      R5,(R0+R2)     R5 <-- 0xF00F000F
        62 => "111010" & "00110" & "00010" & "00000" & "00000010000", -- LWI     R6,16(R2)      R6 <-- 0x7FFFF00F
        64 => "101000" & "00111" & "00000" & "00000" & "00100011000", -- ORI     R7,#280        R7 <-- 280
        65 => "100111" & "00100" & "00000" & "00111" & "00000000000", -- BGT     R0,R7          PC <-- PC + 4
        66 => "100110" & "00000" & "01000" & "00111" & "00000000000", -- BRA     RB             PC <-- 70x4
        ---------------------------------------------------------------------------------------------------------------------------
        70 => "001000" & "00001" & "00000" & "00000" & "00000000001", -- ADDI    R1,R0,#1       R1 <-- 1
        71 => "011001" & "00010" & "00001" & "00000" & "10000000001", -- BSLLI   R2,R1,#1       R2 <-- 2
        72 => "011001" & "00011" & "00010" & "00000" & "11000000010", -- BSLAI   R3,R2,#2       R3 <-- 8
        73 => "011001" & "00100" & "00011" & "00000" & "11000011100", -- BSLLI   R4,R3,#16      R4 <-- 0x80000000
        74 => "011001" & "00101" & "00100" & "00000" & "01000011100", -- BSRAI   R5,R4,#16      R5 <-- 0xFFFFFFF8
        75 => "011001" & "00110" & "00101" & "00000" & "00000000001", -- BSRLI   R6,R5,#1       R6 <-- 0x7FFFFFFC
        76 => "011001" & "00111" & "00110" & "00000" & "01000011100", -- BSRAI   R5,R4,#16      R7 <-- 7
        77 => "101111" & "00001" & "00001" & "00000" & "00000000000", -- BNEI    R1,#0          PC <-- 77x4
        others => x"00000000" -- NOP
);

shared variable RAM : MEM_TYPE := InitValue0;

begin

-----------------------------------------
-- PORT A (read-only)
-----------------------------------------
uRead: process (CLK)
begin
    if rising_edge(CLK) then
        DO_A <= RAM(conv_integer(Addr_A(PC_WIDTH-1 downto 2)));
    end if;
end process;

-----------------------------------------
-- PORT B
-----------------------------------------
process (CLK)
begin
    if rising_edge(CLK) then
        if WE_B='1' then
            RAM(conv_integer(Addr_B(PC_WIDTH-1 downto 2))) := DI_B;
        end if;
        DO_B <= RAM(conv_integer(Addr_B(PC_WIDTH-1 downto 2)));
    end if;
end process;
         
end Behavioral;
